// RISCVmulti.sv
// risc-v multicycle processor
// Christian Johnson
// chrjohnson@hmc.edu
// 12/3/2024

// top module
module top(input  logic        clk, reset,
           output logic [31:0] WriteData, DataAdr,
           output logic        MemWrite);



endmodule

// unified memory module
//      combines both the dmem and imem module from the RISCVsingle processor


// RISCVmulti module containing calls to the controller and datapath modules


// multicycle controller module

//// Main Decoder module
    

//// ALU Decoder module


// Datapath module


// Extend module


// Register File module


// flopr module


// Multiplexers


// 2x1 Mux module


// 3x1 Mux module


// ALU module
